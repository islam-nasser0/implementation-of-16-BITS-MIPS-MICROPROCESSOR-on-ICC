module VCCKHA( inout  VCC);  
endmodule

module GNDKHA( inout  GND);  
endmodule

module VCC3IHA( inout  VCC3I);  
endmodule

module GND3IHA( inout  GND3I);  
endmodule

module CORNERHA( );  
endmodule
